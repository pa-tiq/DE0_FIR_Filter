-- Generic 256 point DIF FFT algorithm using a register
-- array for data and coefficients

--PACKAGE n_bits_int IS          -- User defined types
--	SUBTYPE U9 IS INTEGER RANGE 0 TO 2**9-1;
--	SUBTYPE S16 IS INTEGER RANGE -2**15 TO 2**15-1;
--	SUBTYPE S32 IS INTEGER RANGE -2147483647 TO 2147483647;
--	TYPE ARRAY0_7S16 IS ARRAY (0 TO 7) of S16;
--	TYPE ARRAY0_255S16 IS ARRAY (0 TO 255) of S16;
--	TYPE ARRAY0_127S16 IS ARRAY (0 TO 127) of S16;
--	TYPE STATE_TYPE IS(start, load, calc, update, reverse, done);
--END n_bits_int;

--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
--
--PACKAGE n_bits_int IS          -- User defined types
--	SUBTYPE U9 IS INTEGER RANGE 0 TO 2**9-1;
--	SUBTYPE S16N IS INTEGER RANGE -2**15 TO 2**15-1;
--	SUBTYPE S16 IS STD_LOGIC_VECTOR(15 downto 0);
--	SUBTYPE S16S IS SIGNED(15 downto 0);
--	TYPE ARRAY0_7S16 IS ARRAY (0 TO 7) of S16;
--	TYPE ARRAY0_255S16 IS ARRAY (0 TO 255) of S16;
--	TYPE ARRAY0_255S16S IS ARRAY (0 TO 255) of S16S;
--	TYPE ARRAY0_255S16N IS ARRAY (0 TO 255) of S16N;
--	TYPE ARRAY0_127S16N IS ARRAY (0 TO 127) of S16N;
--	TYPE ARRAY0_127S16S IS ARRAY (0 TO 127) of S16S;
--	TYPE STATE_TYPE IS(start, load, calc, update, reverse, done);
--END n_bits_int;

LIBRARY work; 
USE work.n_bits_int.ALL;

LIBRARY ieee; 
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_signed.ALL;
-- --------------------------------------------------------
ENTITY fft256 IS   ------> Interface
generic ( 	
	LFilter  		: INTEGER 	;
	Log2LFilter     : INTEGER   ); -- Filter length
PORT (
	clk, reset 			: IN  STD_LOGIC; 	-- Clock and reset
	xr_in, xi_in   		: IN  S16; 		 	-- Real and imag. input
	fft_valid 			: OUT STD_LOGIC; 	-- FFT output is valid
	fftr, ffti 			: OUT S16; 		 	-- Real and imag. output
	rcount_o 			: OUT U9; 			-- Bitreverese index counter
	xr_out, xi_out 		: OUT ARRAY0_7S16; 	-- First 8 reg. files
	stage_o, gcount_o 	: OUT U9; 			-- Stage and group count
	i1_o, i2_o 			: OUT U9; 			-- (Dual) data index
	k1_o, k2_o 			: OUT U9; 			-- Index offset
	w_o, dw_o  			: OUT U9; 			-- Cos/Sin (increment) angle
	wo 					: OUT U9);			-- Decision tree location loop FSM
END fft256;

ARCHITECTURE fpga OF fft256 IS

	SIGNAL s    	: STATE_TYPE; -- State machine variable
	--CONSTANT N 	: U9 := 256; -- Number of points
	--CONSTANT ldN 	: U9 := 8; -- Log_2 number of points
	CONSTANT N 		: U9 := LFilter; -- Number of points
	CONSTANT ldN 	: U9 := Log2LFilter; -- Log_2 number of points

	-- Register array for 16 bit precision:
	SIGNAL xr, xi : ARRAY0_255S16;
	--SIGNAL xr, xi 	: ARRAY0_255S16S;
	SIGNAL w: U9 	:= 0;

	-- sine and cosine coefficient arrays RANGE -16379 to 16384

	-- L=127
	-- CONSTANT cos_rom : ARRAY0_127S16 := (
	-- 	16340,16305,16261,16207,16143,16069,15986,15893,15791,15679,15557,15426,15286,15137,14978,14811,14635,14449,14256,14053,13842,13623,13395,13160,12916,12665,12406,12140,11866,11585,11297,11003,10702,10394,10080,9760,9434,9102,8765,8423,8076,7723,7366,7005,6639,6270,5897,5520,5139,4756,4370,3981,3590,3196,2801,2404,2006,1606,1205,804,402,0,-402,-804,-1205,-1606,-2006,-2404,-2801,-3196,-3590,-3981,-4370,-4756,-5139,-5520,-5897,-6270,-6639,-7005,-7366,-7723,-8076,-8423,-8765,-9102,-9434,-9760,-10080,-10394,-10702,-11003,-11297,-11585,-11866,-12140,-12406,-12665,-12916,-13160,-13395,-13623,-13842,-14053,-14256,-14449,-14635,-14811,-14978,-15137,-15286,-15426,-15557,-15679,-15791,-15893,-15986,-16069,-16143,-16207,-16261,-16305,-16340,-16364,-16379
	-- );
	-- CONSTANT sin_rom : ARRAY0_127S16 := (
	-- 	0,402,804,1205,1606,2006,2404,2801,3196,3590,3981,4370,4756,5139,5520,5897,6270,	6639,7005,7366,7723,8076,8423,8765,9102,9434,9760,10080,	10394,10702,11003,11297,11585,11866,12140,12406,12665,12916,	13160,13395,13623,13842,14053,14256,14449,14635,14811,14978,	15137,15286,15426,15557,15679,15791,15893,15986,16069,16143,	16207,16261,16305,16340,16364,16379,16384,16379,16364,16340,	16305,16261,16207,16143,16069,15986,15893,15791,15679,15557,	15426,15286,15137,14978,14811,14635,14449,14256,14053,13842,	13623,13395,13160,12916,12665,12406,12140,11866,11585,11297,	11003,10702,10394,10080,9760,9434,9102,8765,8423,8076,7723,	7366,7005,6639,6270,5897,5520,5139,4756,4370,3981,3590,3196,	2801,2404,2006,1606,1205,804,402
	-- );

	-- L=512 
	--CONSTANT cos_rom : ARRAY0_127S16 := (
	--	16384,16384,16383,16381,16379,16376,16373,16369,16364,16359,16353,16347,16339,16332,16323,16314,16305,16295,16284,16272,16260,16248,16234,16221,16206,16191,16175,16159,16142,16124,16106,16087,16068,16048,16027,16006,15984,15962,15939,15915,15891,15866,15841,15815,15788,15761,15733,15705,15676,15646,15616,15585,15554,15522,15490,15456,15423,15388,15354,15318,15282,15245,15208,15171,15132,15093,15054,15014,14973,14932,14890,14848,14805,14762,14718,14673,14628,14582,14536,14490,14442,14394,14346,14297,14248,14198,14147,14096,14044,13992,13940,13886,13833,13779,13724,13669,13613,13556,13500,13442,13384,13326,13267,13208,13148,13088,13027,12966,12904,12841,12779,12715,12652,12587,12523,12457,12392,12326,12259,12192,12125,12057,11988,11919,11850,11780,11710,11639,11568,11497,11425,11352,11279,11206,11132,11058,10984,10909,10834,10758,10682,10605,10528,10451,10373,10295,10216,10137,10058,9978,9898,9818,9737,9656,9574,9492,9410,9327,9244,9161,9077,8993,8909,8824,8739,8654,8568,8482,8396,8309,8222,8135,8047,7960,7871,7783,7694,7605,7516,7426,7336,7246,7156,7065,6974,6882,6791,6699,6607,6515,6422,6330,6237,6143,6050,5956,5862,5768,5674,5579,5484,5389,5294,5199,5103,5007,4911,4815,4719,4622,4525,4429,4331,4234,4137,4039,3942,3844,3746,3648,3549,3451,3353,3254,3155,3056,2957,2858,2759,2660,2560,2461,2361,2261,2162,2062,1962,1862,1762,1661,1561,1461,1361,1260,1160,1059,959,858,758,657,556,456,355,254,154,53,-48,-149,-249,-350,-451,-551,-652,-753,-853,-954,-1054,-1155,-1255,-1356,-1456,-1556,-1656,-1757,-1857,-1957,-2057,-2157,-2256,-2356,-2456,-2555,-2655,-2754,-2853,-2952,-3051,-3150,-3249,-3348,-3446,-3544,-3643,-3741,-3839,-3937,-4034,-4132,-4229,-4326,-4424,-4520,-4617,-4714,-4810,-4906,-5002,-5098,-5194,-5289,-5384,-5479,-5574,-5669,-5763,-5857,-5951,-6045,-6138,-6232,-6325,-6417,-6510,-6602,-6694,-6786,-6877,-6969,-7060,-7151,-7241,-7331,-7421,-7511,-7600,-7689,-7778,-7866,-7955,-8042,-8130,-8217,-8304,-8391,-8477,-8563,-8649,-8734,-8819,-8904,-8988,-9072,-9156,-9239,-9322,-9405,-9487,-9569,-9651,-9732,-9813,-9893,-9973,-10053,-10132,-10211,-10290,-10368,-10446,-10523,-10600,-10677,-10753,-10829,-10904,-10979,-11053,-11127,-11201,-11274,-11347,-11420,-11492,-11563,-11634,-11705,-11775,-11845,-11914,-11983,-12052,-12120,-12187,-12254,-12321,-12387,-12452,-12518,-12582,-12647,-12710,-12774,-12836,-12899,-12961,-13022,-13083,-13143,-13203,-13262,-13321,-13379,-13437,-13495,-13551,-13608,-13664,-13719,-13774,-13828,-13881,-13935,-13987,-14039,-14091,-14142,-14193,-14243,-14292,-14341,-14389,-14437,-14485,-14531,-14577,-14623,-14668,-14713,-14757,-14800,-14843,-14885,-14927,-14968,-15009,-15049,-15088,-15127,-15166,-15203,-15240,-15277,-15313,-15349,-15383,-15418,-15451,-15485,-15517,-15549,-15580,-15611,-15641,-15671,-15700,-15728,-15756,-15783,-15810,-15836,-15861,-15886,-15910,-15934,-15957,-15979,-16001,-16022,-16043,-16063,-16082,-16101,-16119,-16137,-16154,-16170,-16186,-16201,-16216,-16229,-16243,-16255,-16267,-16279,-16290,-16300,-16309,-16318,-16327,-16334,-16342,-16348,-16354,-16359,-16364,-16368,-16371,-16374,-16376,-16378,-16379,-16379
	--);
	--CONSTANT sin_rom : ARRAY0_127S16 := (
	--	0,101,201,302,403,504,604,705,806,906,1007,1107,1208,1308,1408,1509,1609,1709,1809,1909,2009,2109,2209,2309,2409,2508,2608,2707,2806,2906,3005,3104,3203,3301,3400,3498,3597,3695,3793,3891,3989,4086,4184,4281,4378,4475,4572,4669,4765,4861,4957,5053,5149,5245,5340,5435,5530,5625,5719,5813,5908,6001,6095,6188,6282,6374,6467,6560,6652,6744,6835,6927,7018,7109,7199,7290,7380,7470,7559,7648,7737,7826,7914,8002,8090,8177,8265,8351,8438,8524,8610,8696,8781,8866,8950,9034,9118,9202,9285,9368,9450,9532,9614,9695,9776,9857,9937,10017,10097,10176,10255,10333,10411,10489,10566,10643,10719,10795,10870,10946,11020,11095,11169,11242,11315,11388,11460,11532,11603,11674,11744,11814,11884,11953,12022,12090,12158,12225,12292,12358,12424,12490,12555,12619,12683,12747,12810,12872,12934,12996,13057,13118,13178,13237,13296,13355,13413,13471,13528,13584,13640,13696,13751,13805,13859,13913,13966,14018,14070,14121,14172,14222,14272,14321,14370,14418,14466,14513,14559,14605,14651,14695,14740,14783,14826,14869,14911,14953,14993,15034,15074,15113,15151,15189,15227,15264,15300,15336,15371,15406,15440,15473,15506,15538,15570,15601,15631,15661,15690,15719,15747,15775,15802,15828,15854,15879,15903,15927,15951,15973,15995,16017,16038,16058,16078,16097,16115,16133,16150,16167,16183,16199,16213,16228,16241,16254,16266,16278,16289,16300,16310,16319,16328,16336,16343,16350,16356,16362,16367,16371,16375,16378,16380,16382,16383,16384,16384,16383,16382,16380,16378,16375,16371,16367,16362,16356,16350,16343,16336,16328,16319,16310,16300,16289,16278,16266,16254,16241,16228,16213,16199,16183,16167,16150,16133,16115,16097,16078,16058,16038,16017,15995,15973,15951,15927,15903,15879,15854,15828,15802,15775,15747,15719,15690,15661,15631,15601,15570,15538,15506,15473,15440,15406,15371,15336,15300,15264,15227,15189,15151,15113,15074,15034,14993,14953,14911,14869,14826,14783,14740,14695,14651,14605,14559,14513,14466,14418,14370,14321,14272,14222,14172,14121,14070,14018,13966,13913,13859,13805,13751,13696,13640,13584,13528,13471,13413,13355,13296,13237,13178,13118,13057,12996,12934,12872,12810,12747,12683,12619,12555,12490,12424,12358,12292,12225,12158,12090,12022,11953,11884,11814,11744,11674,11603,11532,11460,11388,11315,11242,11169,11095,11020,10946,10870,10795,10719,10643,10566,10489,10411,10333,10255,10176,10097,10017,9937,9857,9776,9695,9614,9532,9450,9368,9285,9202,9118,9034,8950,8866,8781,8696,8610,8524,8438,8351,8265,8177,8090,8002,7914,7826,7737,7648,7559,7470,7380,7290,7199,7109,7018,6927,6835,6744,6652,6560,6467,6374,6282,6188,6095,6001,5908,5813,5719,5625,5530,5435,5340,5245,5149,5053,4957,4861,4765,4669,4572,4475,4378,4281,4184,4086,3989,3891,3793,3695,3597,3498,3400,3301,3203,3104,3005,2906,2806,2707,2608,2508,2409,2309,2209,2109,2009,1909,1809,1709,1609,1509,1408,1308,1208,1107,1007,906,806,705,604,504,403,302,201,101,0
	--);

	-- L=1024 
	--CONSTANT cos_rom : ARRAY0_127S16 := (
	--	16384,16384,16384,16383,16383,16382,16381,16380,16379,16378,16376,16375,16373,16371,16369,16367,16364,16362,16359,16356,16353,16350,16347,16343,16340,16336,16332,16328,16323,16319,16315,16310,16305,16300,16295,16289,16284,16278,16273,16267,16261,16254,16248,16241,16235,16228,16221,16214,16206,16199,16191,16183,16176,16167,16159,16151,16142,16134,16125,16116,16107,16097,16088,16078,16069,16059,16049,16038,16028,16018,16007,15996,15985,15974,15963,15951,15940,15928,15916,15904,15892,15880,15867,15855,15842,15829,15816,15803,15789,15776,15762,15748,15735,15720,15706,15692,15677,15663,15648,15633,15618,15602,15587,15571,15556,15540,15524,15508,15491,15475,15458,15441,15425,15408,15390,15373,15356,15338,15320,15302,15284,15266,15248,15229,15211,15192,15173,15154,15135,15115,15096,15076,15056,15036,15016,14996,14976,14955,14935,14914,14893,14872,14851,14830,14808,14787,14765,14743,14721,14699,14676,14654,14631,14609,14586,14563,14540,14517,14493,14470,14446,14422,14398,14374,14350,14326,14301,14277,14252,14227,14202,14177,14151,14126,14100,14075,14049,14023,13997,13971,13944,13918,13891,13865,13838,13811,13783,13756,13729,13701,13674,13646,13618,13590,13562,13533,13505,13477,13448,13419,13390,13361,13332,13303,13273,13244,13214,13184,13154,13124,13094,13064,13033,13003,12972,12941,12910,12879,12848,12817,12785,12754,12722,12690,12659,12627,12594,12562,12530,12497,12465,12432,12399,12366,12333,12300,12267,12233,12200,12166,12132,12099,12065,12031,11996,11962,11928,11893,11858,11824,11789,11754,11719,11683,11648,11613,11577,11541,11506,11470,11434,11398,11362,11325,11289,11252,11216,11179,11142,11105,11068,11031,10994,10956,10919,10881,10844,10806,10768,10730,10692,10654,10616,10577,10539,10500,10462,10423,10384,10345,10306,10267,10227,10188,10149,10109,10069,10030,9990,9950,9910,9870,9830,9789,9749,9708,9668,9627,9586,9546,9505,9464,9423,9381,9340,9299,9257,9216,9174,9132,9090,9049,9007,8965,8922,8880,8838,8795,8753,8710,8668,8625,8582,8539,8496,8453,8410,8367,8324,8280,8237,8193,8150,8106,8062,8018,7974,7930,7886,7842,7798,7754,7709,7665,7621,7576,7531,7487,7442,7397,7352,7307,7262,7217,7172,7126,7081,7036,6990,6945,6899,6853,6808,6762,6716,6670,6624,6578,6532,6486,6440,6393,6347,6300,6254,6207,6161,6114,6068,6021,5974,5927,5880,5833,5786,5739,5692,5645,5597,5550,5503,5455,5408,5360,5313,5265,5218,5170,5122,5074,5026,4978,4931,4883,4834,4786,4738,4690,4642,4594,4545,4497,4448,4400,4352,4303,4254,4206,4157,4109,4060,4011,3962,3913,3865,3816,3767,3718,3669,3620,3571,3521,3472,3423,3374,3325,3275,3226,3177,3127,3078,3029,2979,2930,2880,2831,2781,2731,2682,2632,2583,2533,2483,2433,2384,2334,2284,2234,2184,2134,2085,2035,1985,1935,1885,1835,1785,1735,1685,1635,1585,1535,1485,1434,1384,1334,1284,1234,1184,1134,1083,1033,983,933,882,832,782,732,681,631,581,531,480,430,380,329,279,229,179,128,78,28,-23,-73,-123,-174,-224,-274,-324,-375,-425,-475,-526,-576,-626,-676,-727,-777,-827,-877,-928,-978,-1028,-1078,-1129,-1179,-1229,-1279,-1329,-1379,-1429,-1480,-1530,-1580,-1630,-1680,-1730,-1780,-1830,-1880,-1930,-1980,-2030,-2080,-2129,-2179,-2229,-2279,-2329,-2379,-2428,-2478,-2528,-2578,-2627,-2677,-2726,-2776,-2826,-2875,-2925,-2974,-3024,-3073,-3122,-3172,-3221,-3270,-3320,-3369,-3418,-3467,-3516,-3566,-3615,-3664,-3713,-3762,-3811,-3860,-3908,-3957,-4006,-4055,-4104,-4152,-4201,-4249,-4298,-4347,-4395,-4443,-4492,-4540,-4589,-4637,-4685,-4733,-4781,-4829,-4878,-4926,-4973,-5021,-5069,-5117,-5165,-5213,-5260,-5308,-5355,-5403,-5450,-5498,-5545,-5592,-5640,-5687,-5734,-5781,-5828,-5875,-5922,-5969,-6016,-6063,-6109,-6156,-6202,-6249,-6295,-6342,-6388,-6435,-6481,-6527,-6573,-6619,-6665,-6711,-6757,-6803,-6848,-6894,-6940,-6985,-7031,-7076,-7121,-7167,-7212,-7257,-7302,-7347,-7392,-7437,-7482,-7526,-7571,-7616,-7660,-7704,-7749,-7793,-7837,-7881,-7925,-7969,-8013,-8057,-8101,-8145,-8188,-8232,-8275,-8319,-8362,-8405,-8448,-8491,-8534,-8577,-8620,-8663,-8705,-8748,-8790,-8833,-8875,-8917,-8960,-9002,-9044,-9085,-9127,-9169,-9211,-9252,-9294,-9335,-9376,-9418,-9459,-9500,-9541,-9581,-9622,-9663,-9703,-9744,-9784,-9825,-9865,-9905,-9945,-9985,-10025,-10064,-10104,-10144,-10183,-10222,-10262,-10301,-10340,-10379,-10418,-10457,-10495,-10534,-10572,-10611,-10649,-10687,-10725,-10763,-10801,-10839,-10876,-10914,-10951,-10989,-11026,-11063,-11100,-11137,-11174,-11211,-11247,-11284,-11320,-11357,-11393,-11429,-11465,-11501,-11536,-11572,-11608,-11643,-11678,-11714,-11749,-11784,-11819,-11853,-11888,-11923,-11957,-11991,-12026,-12060,-12094,-12127,-12161,-12195,-12228,-12262,-12295,-12328,-12361,-12394,-12427,-12460,-12492,-12525,-12557,-12589,-12622,-12654,-12685,-12717,-12749,-12780,-12812,-12843,-12874,-12905,-12936,-12967,-12998,-13028,-13059,-13089,-13119,-13149,-13179,-13209,-13239,-13268,-13298,-13327,-13356,-13385,-13414,-13443,-13472,-13500,-13528,-13557,-13585,-13613,-13641,-13669,-13696,-13724,-13751,-13778,-13806,-13833,-13860,-13886,-13913,-13939,-13966,-13992,-14018,-14044,-14070,-14095,-14121,-14146,-14172,-14197,-14222,-14247,-14272,-14296,-14321,-14345,-14369,-14393,-14417,-14441,-14465,-14488,-14512,-14535,-14558,-14581,-14604,-14626,-14649,-14671,-14694,-14716,-14738,-14760,-14782,-14803,-14825,-14846,-14867,-14888,-14909,-14930,-14950,-14971,-14991,-15011,-15031,-15051,-15071,-15091,-15110,-15130,-15149,-15168,-15187,-15206,-15224,-15243,-15261,-15279,-15297,-15315,-15333,-15351,-15368,-15385,-15403,-15420,-15436,-15453,-15470,-15486,-15503,-15519,-15535,-15551,-15566,-15582,-15597,-15613,-15628,-15643,-15658,-15672,-15687,-15701,-15715,-15730,-15743,-15757,-15771,-15784,-15798,-15811,-15824,-15837,-15850,-15862,-15875,-15887,-15899,-15911,-15923,-15935,-15946,-15958,-15969,-15980,-15991,-16002,-16013,-16023,-16033,-16044,-16054,-16064,-16073,-16083,-16092,-16102,-16111,-16120,-16129,-16137,-16146,-16154,-16162,-16171,-16178,-16186,-16194,-16201,-16209,-16216,-16223,-16230,-16236,-16243,-16249,-16256,-16262,-16268,-16273,-16279,-16284,-16290,-16295,-16300,-16305,-16310,-16314,-16318,-16323,-16327,-16331,-16335,-16338,-16342,-16345,-16348,-16351,-16354,-16357,-16359,-16362,-16364,-16366,-16368,-16370,-16371,-16373,-16374,-16375,-16376,-16377,-16378,-16378,-16379,-16379,-16379
	--);
	--CONSTANT sin_rom : ARRAY0_127S16 := (
	--	0,50,101,151,201,252,302,352,402,453,503,553,604,654,704,754,805,855,905,955,1006,1056,1106,1156,1206,1257,1307,1357,1407,1457,1507,1557,1607,1658,1708,1758,1808,1858,1908,1958,2008,2057,2107,2157,2207,2257,2307,2357,2406,2456,2506,2556,2605,2655,2705,2754,2804,2853,2903,2952,3002,3051,3101,3150,3199,3249,3298,3347,3397,3446,3495,3544,3593,3642,3691,3740,3789,3838,3887,3936,3985,4034,4082,4131,4180,4228,4277,4325,4374,4422,4471,4519,4568,4616,4664,4712,4761,4809,4857,4905,4953,5001,5049,5096,5144,5192,5240,5287,5335,5382,5430,5477,5525,5572,5619,5667,5714,5761,5808,5855,5902,5949,5996,6043,6089,6136,6183,6229,6276,6322,6369,6415,6461,6507,6553,6600,6646,6692,6737,6783,6829,6875,6920,6966,7011,7057,7102,7148,7193,7238,7283,7328,7373,7418,7463,7508,7552,7597,7641,7686,7730,7775,7819,7863,7907,7951,7995,8039,8083,8127,8170,8214,8257,8301,8344,8387,8430,8474,8517,8560,8602,8645,8688,8731,8773,8816,8858,8900,8942,8984,9027,9068,9110,9152,9194,9235,9277,9318,9360,9401,9442,9483,9524,9565,9606,9647,9687,9728,9768,9809,9849,9889,9929,9969,10009,10049,10088,10128,10167,10207,10246,10285,10324,10363,10402,10441,10480,10519,10557,10596,10634,10672,10710,10748,10786,10824,10862,10899,10937,10974,11012,11049,11086,11123,11160,11197,11233,11270,11306,11343,11379,11415,11451,11487,11523,11559,11594,11630,11665,11700,11735,11771,11805,11840,11875,11910,11944,11979,12013,12047,12081,12115,12149,12182,12216,12249,12283,12316,12349,12382,12415,12448,12481,12513,12545,12578,12610,12642,12674,12706,12738,12769,12801,12832,12863,12894,12925,12956,12987,13017,13048,13078,13109,13139,13169,13199,13228,13258,13287,13317,13346,13375,13404,13433,13462,13490,13519,13547,13575,13604,13632,13659,13687,13715,13742,13769,13797,13824,13851,13878,13904,13931,13957,13983,14010,14036,14062,14087,14113,14138,14164,14189,14214,14239,14264,14289,14313,14338,14362,14386,14410,14434,14458,14481,14505,14528,14551,14574,14597,14620,14643,14665,14687,14710,14732,14754,14775,14797,14819,14840,14861,14882,14903,14924,14945,14965,14986,15006,15026,15046,15066,15086,15105,15125,15144,15163,15182,15201,15220,15238,15257,15275,15293,15311,15329,15347,15364,15382,15399,15416,15433,15450,15466,15483,15499,15516,15532,15548,15563,15579,15595,15610,15625,15640,15655,15670,15684,15699,15713,15727,15741,15755,15769,15783,15796,15809,15822,15835,15848,15861,15874,15886,15898,15910,15922,15934,15946,15957,15968,15980,15991,16002,16012,16023,16033,16044,16054,16064,16073,16083,16093,16102,16111,16120,16129,16138,16147,16155,16163,16172,16180,16187,16195,16203,16210,16217,16224,16231,16238,16245,16251,16257,16264,16270,16275,16281,16287,16292,16297,16302,16307,16312,16317,16321,16326,16330,16334,16338,16341,16345,16348,16352,16355,16358,16360,16363,16365,16368,16370,16372,16374,16376,16377,16378,16380,16381,16382,16382,16383,16384,16384,16384,16384,16384,16384,16383,16382,16382,16381,16380,16378,16377,16376,16374,16372,16370,16368,16365,16363,16360,16358,16355,16352,16348,16345,16341,16338,16334,16330,16326,16321,16317,16312,16307,16302,16297,16292,16287,16281,16275,16270,16264,16257,16251,16245,16238,16231,16224,16217,16210,16203,16195,16187,16180,16172,16163,16155,16147,16138,16129,16120,16111,16102,16093,16083,16073,16064,16054,16044,16033,16023,16012,16002,15991,15980,15968,15957,15946,15934,15922,15910,15898,15886,15874,15861,15848,15835,15822,15809,15796,15783,15769,15755,15741,15727,15713,15699,15684,15670,15655,15640,15625,15610,15595,15579,15563,15548,15532,15516,15499,15483,15466,15450,15433,15416,15399,15382,15364,15347,15329,15311,15293,15275,15257,15238,15220,15201,15182,15163,15144,15125,15105,15086,15066,15046,15026,15006,14986,14965,14945,14924,14903,14882,14861,14840,14819,14797,14775,14754,14732,14710,14687,14665,14643,14620,14597,14574,14551,14528,14505,14481,14458,14434,14410,14386,14362,14338,14313,14289,14264,14239,14214,14189,14164,14138,14113,14087,14062,14036,14010,13983,13957,13931,13904,13878,13851,13824,13797,13769,13742,13715,13687,13659,13632,13604,13575,13547,13519,13490,13462,13433,13404,13375,13346,13317,13287,13258,13228,13199,13169,13139,13109,13078,13048,13017,12987,12956,12925,12894,12863,12832,12801,12769,12738,12706,12674,12642,12610,12578,12545,12513,12481,12448,12415,12382,12349,12316,12283,12249,12216,12182,12149,12115,12081,12047,12013,11979,11944,11910,11875,11840,11805,11771,11735,11700,11665,11630,11594,11559,11523,11487,11451,11415,11379,11343,11306,11270,11233,11197,11160,11123,11086,11049,11012,10974,10937,10899,10862,10824,10786,10748,10710,10672,10634,10596,10557,10519,10480,10441,10402,10363,10324,10285,10246,10207,10167,10128,10088,10049,10009,9969,9929,9889,9849,9809,9768,9728,9687,9647,9606,9565,9524,9483,9442,9401,9360,9318,9277,9235,9194,9152,9110,9068,9027,8984,8942,8900,8858,8816,8773,8731,8688,8645,8602,8560,8517,8474,8430,8387,8344,8301,8257,8214,8170,8127,8083,8039,7995,7951,7907,7863,7819,7775,7730,7686,7641,7597,7552,7508,7463,7418,7373,7328,7283,7238,7193,7148,7102,7057,7011,6966,6920,6875,6829,6783,6737,6692,6646,6600,6553,6507,6461,6415,6369,6322,6276,6229,6183,6136,6089,6043,5996,5949,5902,5855,5808,5761,5714,5667,5619,5572,5525,5477,5430,5382,5335,5287,5240,5192,5144,5096,5049,5001,4953,4905,4857,4809,4761,4712,4664,4616,4568,4519,4471,4422,4374,4325,4277,4228,4180,4131,4082,4034,3985,3936,3887,3838,3789,3740,3691,3642,3593,3544,3495,3446,3397,3347,3298,3249,3199,3150,3101,3051,3002,2952,2903,2853,2804,2754,2705,2655,2605,2556,2506,2456,2406,2357,2307,2257,2207,2157,2107,2057,2008,1958,1908,1858,1808,1758,1708,1658,1607,1557,1507,1457,1407,1357,1307,1257,1206,1156,1106,1056,1006,955,905,855,805,754,704,654,604,553,503,453,402,352,302,252,201,151,101,50,0
	--);
	
	-- L=2048 
	CONSTANT cos_rom : ARRAY0_127S16 := (
		16384,16384,16384,16384,16384,16384,16383,16383,16383,16382,16382,16382,16381,16381,16380,16380,16379,16378,16378,16377,16376,16375,16375,16374,16373,16372,16371,16370,16369,16368,16367,16365,16364,16363,16362,16360,16359,16358,16356,16355,16353,16352,16350,16348,16347,16345,16343,16341,16340,16338,16336,16334,16332,16330,16328,16326,16324,16321,16319,16317,16315,16312,16310,16307,16305,16303,16300,16297,16295,16292,16290,16287,16284,16281,16278,16276,16273,16270,16267,16264,16261,16258,16254,16251,16248,16245,16242,16238,16235,16231,16228,16224,16221,16217,16214,16210,16207,16203,16199,16195,16191,16188,16184,16180,16176,16172,16168,16164,16159,16155,16151,16147,16143,16138,16134,16130,16125,16121,16116,16112,16107,16102,16098,16093,16088,16083,16079,16074,16069,16064,16059,16054,16049,16044,16039,16034,16028,16023,16018,16013,16007,16002,15997,15991,15986,15980,15974,15969,15963,15958,15952,15946,15940,15934,15929,15923,15917,15911,15905,15899,15893,15886,15880,15874,15868,15862,15855,15849,15842,15836,15830,15823,15817,15810,15803,15797,15790,15783,15777,15770,15763,15756,15749,15742,15735,15728,15721,15714,15707,15700,15692,15685,15678,15671,15663,15656,15648,15641,15633,15626,15618,15611,15603,15595,15588,15580,15572,15564,15556,15548,15541,15533,15525,15516,15508,15500,15492,15484,15476,15467,15459,15451,15442,15434,15425,15417,15408,15400,15391,15383,15374,15365,15357,15348,15339,15330,15321,15312,15303,15294,15285,15276,15267,15258,15249,15240,15230,15221,15212,15202,15193,15184,15174,15165,15155,15145,15136,15126,15117,15107,15097,15087,15077,15068,15058,15048,15038,15028,15018,15008,14998,14987,14977,14967,14957,14947,14936,14926,14915,14905,14895,14884,14874,14863,14852,14842,14831,14820,14810,14799,14788,14777,14766,14755,14745,14734,14723,14711,14700,14689,14678,14667,14656,14644,14633,14622,14610,14599,14588,14576,14565,14553,14542,14530,14518,14507,14495,14483,14471,14460,14448,14436,14424,14412,14400,14388,14376,14364,14352,14340,14328,14315,14303,14291,14279,14266,14254,14241,14229,14216,14204,14191,14179,14166,14154,14141,14128,14115,14103,14090,14077,14064,14051,14038,14025,14012,13999,13986,13973,13960,13947,13933,13920,13907,13894,13880,13867,13853,13840,13827,13813,13800,13786,13772,13759,13745,13731,13718,13704,13690,13676,13662,13648,13635,13621,13607,13593,13579,13564,13550,13536,13522,13508,13494,13479,13465,13451,13436,13422,13407,13393,13378,13364,13349,13335,13320,13305,13291,13276,13261,13247,13232,13217,13202,13187,13172,13157,13142,13127,13112,13097,13082,13067,13052,13036,13021,13006,12991,12975,12960,12944,12929,12914,12898,12883,12867,12851,12836,12820,12804,12789,12773,12757,12741,12726,12710,12694,12678,12662,12646,12630,12614,12598,12582,12566,12550,12533,12517,12501,12485,12468,12452,12436,12419,12403,12387,12370,12354,12337,12320,12304,12287,12271,12254,12237,12221,12204,12187,12170,12153,12136,12120,12103,12086,12069,12052,12035,12018,12000,11983,11966,11949,11932,11914,11897,11880,11863,11845,11828,11810,11793,11775,11758,11740,11723,11705,11688,11670,11652,11635,11617,11599,11582,11564,11546,11528,11510,11492,11474,11456,11438,11420,11402,11384,11366,11348,11330,11312,11294,11275,11257,11239,11220,11202,11184,11165,11147,11129,11110,11092,11073,11054,11036,11017,10999,10980,10961,10943,10924,10905,10886,10868,10849,10830,10811,10792,10773,10754,10735,10716,10697,10678,10659,10640,10621,10602,10583,10563,10544,10525,10506,10486,10467,10448,10428,10409,10389,10370,10350,10331,10311,10292,10272,10253,10233,10213,10194,10174,10154,10135,10115,10095,10075,10055,10035,10016,9996,9976,9956,9936,9916,9896,9876,9856,9836,9815,9795,9775,9755,9735,9715,9694,9674,9654,9633,9613,9593,9572,9552,9531,9511,9490,9470,9449,9429,9408,9388,9367,9346,9326,9305,9284,9264,9243,9222,9201,9181,9160,9139,9118,9097,9076,9055,9034,9013,8992,8971,8950,8929,8908,8887,8866,8845,8823,8802,8781,8760,8739,8717,8696,8675,8653,8632,8611,8589,8568,8546,8525,8503,8482,8460,8439,8417,8396,8374,8352,8331,8309,8287,8266,8244,8222,8201,8179,8157,8135,8113,8091,8070,8048,8026,8004,7982,7960,7938,7916,7894,7872,7850,7828,7806,7784,7761,7739,7717,7695,7673,7650,7628,7606,7584,7561,7539,7517,7494,7472,7450,7427,7405,7382,7360,7337,7315,7292,7270,7247,7225,7202,7180,7157,7134,7112,7089,7066,7044,7021,6998,6976,6953,6930,6907,6884,6862,6839,6816,6793,6770,6747,6724,6701,6678,6656,6633,6610,6587,6563,6540,6517,6494,6471,6448,6425,6402,6379,6356,6332,6309,6286,6263,6239,6216,6193,6170,6146,6123,6100,6076,6053,6030,6006,5983,5959,5936,5913,5889,5866,5842,5819,5795,5772,5748,5725,5701,5677,5654,5630,5607,5583,5559,5536,5512,5488,5465,5441,5417,5393,5370,5346,5322,5298,5275,5251,5227,5203,5179,5155,5132,5108,5084,5060,5036,5012,4988,4964,4940,4916,4892,4868,4844,4820,4796,4772,4748,4724,4700,4676,4652,4628,4603,4579,4555,4531,4507,4483,4458,4434,4410,4386,4362,4337,4313,4289,4265,4240,4216,4192,4167,4143,4119,4094,4070,4046,4021,3997,3973,3948,3924,3899,3875,3851,3826,3802,3777,3753,3728,3704,3679,3655,3630,3606,3581,3557,3532,3508,3483,3458,3434,3409,3385,3360,3335,3311,3286,3262,3237,3212,3188,3163,3138,3114,3089,3064,3039,3015,2990,2965,2941,2916,2891,2866,2842,2817,2792,2767,2743,2718,2693,2668,2643,2619,2594,2569,2544,2519,2494,2469,2445,2420,2395,2370,2345,2320,2295,2270,2246,2221,2196,2171,2146,2121,2096,2071,2046,2021,1996,1971,1946,1921,1896,1871,1846,1821,1796,1771,1747,1722,1696,1671,1646,1621,1596,1571,1546,1521,1496,1471,1446,1421,1396,1371,1346,1321,1296,1271,1246,1221,1196,1171,1145,1120,1095,1070,1045,1020,995,970,945,920,895,869,844,819,794,769,744,719,694,669,643,618,593,568,543,518,493,468,442,417,392,367,342,317,292,266,241,216,191,166,141,116,90,65,40,15,-10,-35,-60,-85,-111,-136,-161,-186,-211,-236,-261,-287,-312,-337,-362,-387,-412,-437,-463,-488,-513,-538,-563,-588,-613,-638,-664,-689,-714,-739,-764,-789,-814,-839,-864,-890,-915,-940,-965,-990,-1015,-1040,-1065,-1090,-1115,-1140,-1166,-1191,-1216,-1241,-1266,-1291,-1316,-1341,-1366,-1391,-1416,-1441,-1466,-1491,-1516,-1541,-1566,-1591,-1616,-1641,-1666,-1691,-1717,-1742,-1766,-1791,-1816,-1841,-1866,-1891,-1916,-1941,-1966,-1991,-2016,-2041,-2066,-2091,-2116,-2141,-2166,-2191,-2216,-2241,-2265,-2290,-2315,-2340,-2365,-2390,-2415,-2440,-2464,-2489,-2514,-2539,-2564,-2589,-2614,-2638,-2663,-2688,-2713,-2738,-2762,-2787,-2812,-2837,-2861,-2886,-2911,-2936,-2960,-2985,-3010,-3034,-3059,-3084,-3109,-3133,-3158,-3183,-3207,-3232,-3257,-3281,-3306,-3330,-3355,-3380,-3404,-3429,-3453,-3478,-3503,-3527,-3552,-3576,-3601,-3625,-3650,-3674,-3699,-3723,-3748,-3772,-3797,-3821,-3846,-3870,-3894,-3919,-3943,-3968,-3992,-4016,-4041,-4065,-4089,-4114,-4138,-4162,-4187,-4211,-4235,-4260,-4284,-4308,-4332,-4357,-4381,-4405,-4429,-4453,-4478,-4502,-4526,-4550,-4574,-4598,-4623,-4647,-4671,-4695,-4719,-4743,-4767,-4791,-4815,-4839,-4863,-4887,-4911,-4935,-4959,-4983,-5007,-5031,-5055,-5079,-5103,-5127,-5150,-5174,-5198,-5222,-5246,-5270,-5293,-5317,-5341,-5365,-5388,-5412,-5436,-5460,-5483,-5507,-5531,-5554,-5578,-5602,-5625,-5649,-5672,-5696,-5720,-5743,-5767,-5790,-5814,-5837,-5861,-5884,-5908,-5931,-5954,-5978,-6001,-6025,-6048,-6071,-6095,-6118,-6141,-6165,-6188,-6211,-6234,-6258,-6281,-6304,-6327,-6351,-6374,-6397,-6420,-6443,-6466,-6489,-6512,-6535,-6558,-6582,-6605,-6628,-6651,-6673,-6696,-6719,-6742,-6765,-6788,-6811,-6834,-6857,-6879,-6902,-6925,-6948,-6971,-6993,-7016,-7039,-7061,-7084,-7107,-7129,-7152,-7175,-7197,-7220,-7242,-7265,-7287,-7310,-7332,-7355,-7377,-7400,-7422,-7445,-7467,-7489,-7512,-7534,-7556,-7579,-7601,-7623,-7645,-7668,-7690,-7712,-7734,-7756,-7779,-7801,-7823,-7845,-7867,-7889,-7911,-7933,-7955,-7977,-7999,-8021,-8043,-8065,-8086,-8108,-8130,-8152,-8174,-8196,-8217,-8239,-8261,-8282,-8304,-8326,-8347,-8369,-8391,-8412,-8434,-8455,-8477,-8498,-8520,-8541,-8563,-8584,-8606,-8627,-8648,-8670,-8691,-8712,-8734,-8755,-8776,-8797,-8818,-8840,-8861,-8882,-8903,-8924,-8945,-8966,-8987,-9008,-9029,-9050,-9071,-9092,-9113,-9134,-9155,-9176,-9196,-9217,-9238,-9259,-9279,-9300,-9321,-9341,-9362,-9383,-9403,-9424,-9444,-9465,-9485,-9506,-9526,-9547,-9567,-9588,-9608,-9628,-9649,-9669,-9689,-9710,-9730,-9750,-9770,-9790,-9810,-9831,-9851,-9871,-9891,-9911,-9931,-9951,-9971,-9991,-10011,-10030,-10050,-10070,-10090,-10110,-10130,-10149,-10169,-10189,-10208,-10228,-10248,-10267,-10287,-10306,-10326,-10345,-10365,-10384,-10404,-10423,-10443,-10462,-10481,-10501,-10520,-10539,-10558,-10578,-10597,-10616,-10635,-10654,-10673,-10692,-10711,-10730,-10749,-10768,-10787,-10806,-10825,-10844,-10863,-10881,-10900,-10919,-10938,-10956,-10975,-10994,-11012,-11031,-11049,-11068,-11087,-11105,-11124,-11142,-11160,-11179,-11197,-11215,-11234,-11252,-11270,-11289,-11307,-11325,-11343,-11361,-11379,-11397,-11415,-11433,-11451,-11469,-11487,-11505,-11523,-11541,-11559,-11577,-11594,-11612,-11630,-11647,-11665,-11683,-11700,-11718,-11735,-11753,-11770,-11788,-11805,-11823,-11840,-11858,-11875,-11892,-11909,-11927,-11944,-11961,-11978,-11995,-12013,-12030,-12047,-12064,-12081,-12098,-12115,-12131,-12148,-12165,-12182,-12199,-12216,-12232,-12249,-12266,-12282,-12299,-12315,-12332,-12349,-12365,-12382,-12398,-12414,-12431,-12447,-12463,-12480,-12496,-12512,-12528,-12545,-12561,-12577,-12593,-12609,-12625,-12641,-12657,-12673,-12689,-12705,-12721,-12736,-12752,-12768,-12784,-12799,-12815,-12831,-12846,-12862,-12878,-12893,-12909,-12924,-12939,-12955,-12970,-12986,-13001,-13016,-13031,-13047,-13062,-13077,-13092,-13107,-13122,-13137,-13152,-13167,-13182,-13197,-13212,-13227,-13242,-13256,-13271,-13286,-13300,-13315,-13330,-13344,-13359,-13373,-13388,-13402,-13417,-13431,-13446,-13460,-13474,-13489,-13503,-13517,-13531,-13545,-13559,-13574,-13588,-13602,-13616,-13630,-13643,-13657,-13671,-13685,-13699,-13713,-13726,-13740,-13754,-13767,-13781,-13795,-13808,-13822,-13835,-13848,-13862,-13875,-13889,-13902,-13915,-13928,-13942,-13955,-13968,-13981,-13994,-14007,-14020,-14033,-14046,-14059,-14072,-14085,-14098,-14110,-14123,-14136,-14149,-14161,-14174,-14186,-14199,-14211,-14224,-14236,-14249,-14261,-14274,-14286,-14298,-14310,-14323,-14335,-14347,-14359,-14371,-14383,-14395,-14407,-14419,-14431,-14443,-14455,-14466,-14478,-14490,-14502,-14513,-14525,-14537,-14548,-14560,-14571,-14583,-14594,-14605,-14617,-14628,-14639,-14651,-14662,-14673,-14684,-14695,-14706,-14718,-14729,-14740,-14750,-14761,-14772,-14783,-14794,-14805,-14815,-14826,-14837,-14847,-14858,-14869,-14879,-14890,-14900,-14910,-14921,-14931,-14942,-14952,-14962,-14972,-14982,-14993,-15003,-15013,-15023,-15033,-15043,-15053,-15063,-15072,-15082,-15092,-15102,-15112,-15121,-15131,-15140,-15150,-15160,-15169,-15179,-15188,-15197,-15207,-15216,-15225,-15235,-15244,-15253,-15262,-15271,-15280,-15289,-15298,-15307,-15316,-15325,-15334,-15343,-15352,-15360,-15369,-15378,-15386,-15395,-15403,-15412,-15420,-15429,-15437,-15446,-15454,-15462,-15471,-15479,-15487,-15495,-15503,-15511,-15520,-15528,-15536,-15543,-15551,-15559,-15567,-15575,-15583,-15590,-15598,-15606,-15613,-15621,-15628,-15636,-15643,-15651,-15658,-15666,-15673,-15680,-15687,-15695,-15702,-15709,-15716,-15723,-15730,-15737,-15744,-15751,-15758,-15765,-15772,-15778,-15785,-15792,-15798,-15805,-15812,-15818,-15825,-15831,-15837,-15844,-15850,-15857,-15863,-15869,-15875,-15881,-15888,-15894,-15900,-15906,-15912,-15918,-15924,-15929,-15935,-15941,-15947,-15953,-15958,-15964,-15969,-15975,-15981,-15986,-15992,-15997,-16002,-16008,-16013,-16018,-16023,-16029,-16034,-16039,-16044,-16049,-16054,-16059,-16064,-16069,-16074,-16078,-16083,-16088,-16093,-16097,-16102,-16107,-16111,-16116,-16120,-16125,-16129,-16133,-16138,-16142,-16146,-16150,-16154,-16159,-16163,-16167,-16171,-16175,-16179,-16183,-16186,-16190,-16194,-16198,-16202,-16205,-16209,-16212,-16216,-16219,-16223,-16226,-16230,-16233,-16237,-16240,-16243,-16246,-16249,-16253,-16256,-16259,-16262,-16265,-16268,-16271,-16273,-16276,-16279,-16282,-16285,-16287,-16290,-16292,-16295,-16298,-16300,-16302,-16305,-16307,-16310,-16312,-16314,-16316,-16319,-16321,-16323,-16325,-16327,-16329,-16331,-16333,-16335,-16336,-16338,-16340,-16342,-16343,-16345,-16347,-16348,-16350,-16351,-16353,-16354,-16355,-16357,-16358,-16359,-16360,-16362,-16363,-16364,-16365,-16366,-16367,-16368,-16369,-16370,-16370,-16371,-16372,-16373,-16373,-16374,-16375,-16375,-16376,-16376,-16377,-16377,-16377,-16378,-16378,-16378,-16379,-16379,-16379,-16379,-16379,-16379
	);
	CONSTANT sin_rom : ARRAY0_127S16 := (
		0,25,50,75,101,126,151,176,201,226,251,277,302,327,352,377,402,427,453,478,503,528,553,578,603,628,654,679,704,729,754,779,804,829,855,880,905,930,955,980,1005,1030,1055,1080,1106,1131,1156,1181,1206,1231,1256,1281,1306,1331,1356,1381,1406,1431,1456,1482,1507,1532,1557,1582,1607,1632,1657,1682,1707,1732,1757,1782,1807,1832,1857,1882,1907,1932,1957,1982,2007,2032,2056,2081,2106,2131,2156,2181,2206,2231,2256,2281,2306,2331,2355,2380,2405,2430,2455,2480,2505,2529,2554,2579,2604,2629,2654,2678,2703,2728,2753,2778,2802,2827,2852,2877,2901,2926,2951,2976,3000,3025,3050,3075,3099,3124,3149,3173,3198,3223,3247,3272,3296,3321,3346,3370,3395,3420,3444,3469,3493,3518,3542,3567,3591,3616,3641,3665,3690,3714,3739,3763,3787,3812,3836,3861,3885,3910,3934,3958,3983,4007,4032,4056,4080,4105,4129,4153,4178,4202,4226,4251,4275,4299,4323,4348,4372,4396,4420,4445,4469,4493,4517,4541,4565,4590,4614,4638,4662,4686,4710,4734,4758,4782,4806,4830,4854,4878,4902,4926,4950,4974,4998,5022,5046,5070,5094,5118,5142,5166,5190,5213,5237,5261,5285,5309,5332,5356,5380,5404,5427,5451,5475,5499,5522,5546,5570,5593,5617,5640,5664,5688,5711,5735,5758,5782,5805,5829,5852,5876,5899,5923,5946,5970,5993,6016,6040,6063,6086,6110,6133,6156,6180,6203,6226,6250,6273,6296,6319,6342,6366,6389,6412,6435,6458,6481,6504,6527,6550,6574,6597,6620,6643,6666,6688,6711,6734,6757,6780,6803,6826,6849,6872,6894,6917,6940,6963,6986,7008,7031,7054,7076,7099,7122,7144,7167,7190,7212,7235,7257,7280,7302,7325,7347,7370,7392,7415,7437,7459,7482,7504,7527,7549,7571,7593,7616,7638,7660,7682,7705,7727,7749,7771,7793,7815,7837,7860,7882,7904,7926,7948,7970,7992,8014,8035,8057,8079,8101,8123,8145,8167,8188,8210,8232,8254,8275,8297,8319,8340,8362,8384,8405,8427,8448,8470,8491,8513,8534,8556,8577,8599,8620,8641,8663,8684,8705,8727,8748,8769,8790,8812,8833,8854,8875,8896,8917,8938,8960,8981,9002,9023,9044,9065,9085,9106,9127,9148,9169,9190,9211,9231,9252,9273,9294,9314,9335,9356,9376,9397,9417,9438,9459,9479,9500,9520,9541,9561,9581,9602,9622,9642,9663,9683,9703,9724,9744,9764,9784,9804,9825,9845,9865,9885,9905,9925,9945,9965,9985,10005,10025,10044,10064,10084,10104,10124,10143,10163,10183,10203,10222,10242,10262,10281,10301,10320,10340,10359,10379,10398,10418,10437,10456,10476,10495,10514,10534,10553,10572,10591,10610,10630,10649,10668,10687,10706,10725,10744,10763,10782,10801,10820,10839,10857,10876,10895,10914,10932,10951,10970,10989,11007,11026,11044,11063,11081,11100,11118,11137,11155,11174,11192,11210,11229,11247,11265,11284,11302,11320,11338,11356,11374,11393,11411,11429,11447,11465,11483,11500,11518,11536,11554,11572,11590,11607,11625,11643,11661,11678,11696,11713,11731,11749,11766,11784,11801,11818,11836,11853,11871,11888,11905,11922,11940,11957,11974,11991,12008,12025,12042,12059,12076,12093,12110,12127,12144,12161,12178,12195,12212,12228,12245,12262,12278,12295,12312,12328,12345,12361,12378,12394,12411,12427,12443,12460,12476,12492,12509,12525,12541,12557,12573,12589,12605,12622,12638,12654,12669,12685,12701,12717,12733,12749,12765,12780,12796,12812,12827,12843,12859,12874,12890,12905,12921,12936,12952,12967,12982,12998,13013,13028,13043,13059,13074,13089,13104,13119,13134,13149,13164,13179,13194,13209,13224,13239,13253,13268,13283,13298,13312,13327,13342,13356,13371,13385,13400,13414,13429,13443,13457,13472,13486,13500,13514,13529,13543,13557,13571,13585,13599,13613,13627,13641,13655,13669,13683,13697,13710,13724,13738,13752,13765,13779,13792,13806,13819,13833,13846,13860,13873,13887,13900,13913,13926,13940,13953,13966,13979,13992,14005,14018,14031,14044,14057,14070,14083,14096,14109,14121,14134,14147,14160,14172,14185,14197,14210,14222,14235,14247,14260,14272,14284,14297,14309,14321,14333,14346,14358,14370,14382,14394,14406,14418,14430,14442,14453,14465,14477,14489,14501,14512,14524,14536,14547,14559,14570,14582,14593,14605,14616,14627,14639,14650,14661,14672,14683,14695,14706,14717,14728,14739,14750,14761,14772,14782,14793,14804,14815,14826,14836,14847,14858,14868,14879,14889,14900,14910,14920,14931,14941,14951,14962,14972,14982,14992,15002,15013,15023,15033,15043,15053,15062,15072,15082,15092,15102,15111,15121,15131,15140,15150,15160,15169,15179,15188,15197,15207,15216,15225,15235,15244,15253,15262,15271,15281,15290,15299,15308,15317,15325,15334,15343,15352,15361,15369,15378,15387,15395,15404,15413,15421,15430,15438,15446,15455,15463,15471,15480,15488,15496,15504,15512,15520,15528,15536,15544,15552,15560,15568,15576,15584,15591,15599,15607,15614,15622,15630,15637,15645,15652,15659,15667,15674,15681,15689,15696,15703,15710,15717,15725,15732,15739,15746,15752,15759,15766,15773,15780,15787,15793,15800,15807,15813,15820,15826,15833,15839,15846,15852,15858,15865,15871,15877,15883,15889,15896,15902,15908,15914,15920,15926,15931,15937,15943,15949,15955,15960,15966,15972,15977,15983,15988,15994,15999,16005,16010,16015,16021,16026,16031,16036,16041,16046,16051,16056,16061,16066,16071,16076,16081,16086,16091,16095,16100,16105,16109,16114,16118,16123,16127,16132,16136,16140,16145,16149,16153,16157,16162,16166,16170,16174,16178,16182,16186,16190,16193,16197,16201,16205,16208,16212,16216,16219,16223,16226,16230,16233,16236,16240,16243,16246,16250,16253,16256,16259,16262,16265,16268,16271,16274,16277,16280,16283,16285,16288,16291,16294,16296,16299,16301,16304,16306,16309,16311,16313,16316,16318,16320,16322,16325,16327,16329,16331,16333,16335,16337,16339,16340,16342,16344,16346,16348,16349,16351,16352,16354,16355,16357,16358,16360,16361,16362,16364,16365,16366,16367,16368,16369,16370,16371,16372,16373,16374,16375,16376,16377,16377,16378,16379,16379,16380,16380,16381,16381,16382,16382,16383,16383,16383,16383,16384,16384,16384,16384,16384,16384,16384,16384,16384,16384,16383,16383,16383,16383,16382,16382,16381,16381,16380,16380,16379,16379,16378,16377,16377,16376,16375,16374,16373,16372,16371,16370,16369,16368,16367,16366,16365,16364,16362,16361,16360,16358,16357,16355,16354,16352,16351,16349,16348,16346,16344,16342,16340,16339,16337,16335,16333,16331,16329,16327,16325,16322,16320,16318,16316,16313,16311,16309,16306,16304,16301,16299,16296,16294,16291,16288,16285,16283,16280,16277,16274,16271,16268,16265,16262,16259,16256,16253,16250,16246,16243,16240,16236,16233,16230,16226,16223,16219,16216,16212,16208,16205,16201,16197,16193,16190,16186,16182,16178,16174,16170,16166,16162,16157,16153,16149,16145,16140,16136,16132,16127,16123,16118,16114,16109,16105,16100,16095,16091,16086,16081,16076,16071,16066,16061,16056,16051,16046,16041,16036,16031,16026,16021,16015,16010,16005,15999,15994,15988,15983,15977,15972,15966,15960,15955,15949,15943,15937,15931,15926,15920,15914,15908,15902,15896,15889,15883,15877,15871,15865,15858,15852,15846,15839,15833,15826,15820,15813,15807,15800,15793,15787,15780,15773,15766,15759,15752,15746,15739,15732,15725,15717,15710,15703,15696,15689,15681,15674,15667,15659,15652,15645,15637,15630,15622,15614,15607,15599,15591,15584,15576,15568,15560,15552,15544,15536,15528,15520,15512,15504,15496,15488,15480,15471,15463,15455,15446,15438,15430,15421,15413,15404,15395,15387,15378,15369,15361,15352,15343,15334,15325,15317,15308,15299,15290,15281,15271,15262,15253,15244,15235,15225,15216,15207,15197,15188,15179,15169,15160,15150,15140,15131,15121,15111,15102,15092,15082,15072,15062,15053,15043,15033,15023,15013,15002,14992,14982,14972,14962,14951,14941,14931,14920,14910,14900,14889,14879,14868,14858,14847,14836,14826,14815,14804,14793,14782,14772,14761,14750,14739,14728,14717,14706,14695,14683,14672,14661,14650,14639,14627,14616,14605,14593,14582,14570,14559,14547,14536,14524,14512,14501,14489,14477,14465,14453,14442,14430,14418,14406,14394,14382,14370,14358,14346,14333,14321,14309,14297,14284,14272,14260,14247,14235,14222,14210,14197,14185,14172,14160,14147,14134,14121,14109,14096,14083,14070,14057,14044,14031,14018,14005,13992,13979,13966,13953,13940,13926,13913,13900,13887,13873,13860,13846,13833,13819,13806,13792,13779,13765,13752,13738,13724,13710,13697,13683,13669,13655,13641,13627,13613,13599,13585,13571,13557,13543,13529,13514,13500,13486,13472,13457,13443,13429,13414,13400,13385,13371,13356,13342,13327,13312,13298,13283,13268,13253,13239,13224,13209,13194,13179,13164,13149,13134,13119,13104,13089,13074,13059,13043,13028,13013,12998,12982,12967,12952,12936,12921,12905,12890,12874,12859,12843,12827,12812,12796,12780,12765,12749,12733,12717,12701,12685,12669,12654,12638,12622,12605,12589,12573,12557,12541,12525,12509,12492,12476,12460,12443,12427,12411,12394,12378,12361,12345,12328,12312,12295,12278,12262,12245,12228,12212,12195,12178,12161,12144,12127,12110,12093,12076,12059,12042,12025,12008,11991,11974,11957,11940,11922,11905,11888,11871,11853,11836,11818,11801,11784,11766,11749,11731,11713,11696,11678,11661,11643,11625,11607,11590,11572,11554,11536,11518,11500,11483,11465,11447,11429,11411,11393,11374,11356,11338,11320,11302,11284,11265,11247,11229,11210,11192,11174,11155,11137,11118,11100,11081,11063,11044,11026,11007,10989,10970,10951,10932,10914,10895,10876,10857,10839,10820,10801,10782,10763,10744,10725,10706,10687,10668,10649,10630,10610,10591,10572,10553,10534,10514,10495,10476,10456,10437,10418,10398,10379,10359,10340,10320,10301,10281,10262,10242,10222,10203,10183,10163,10143,10124,10104,10084,10064,10044,10025,10005,9985,9965,9945,9925,9905,9885,9865,9845,9825,9804,9784,9764,9744,9724,9703,9683,9663,9642,9622,9602,9581,9561,9541,9520,9500,9479,9459,9438,9417,9397,9376,9356,9335,9314,9294,9273,9252,9231,9211,9190,9169,9148,9127,9106,9085,9065,9044,9023,9002,8981,8960,8938,8917,8896,8875,8854,8833,8812,8790,8769,8748,8727,8705,8684,8663,8641,8620,8599,8577,8556,8534,8513,8491,8470,8448,8427,8405,8384,8362,8340,8319,8297,8275,8254,8232,8210,8188,8167,8145,8123,8101,8079,8057,8035,8014,7992,7970,7948,7926,7904,7882,7860,7837,7815,7793,7771,7749,7727,7705,7682,7660,7638,7616,7593,7571,7549,7527,7504,7482,7459,7437,7415,7392,7370,7347,7325,7302,7280,7257,7235,7212,7190,7167,7144,7122,7099,7076,7054,7031,7008,6986,6963,6940,6917,6894,6872,6849,6826,6803,6780,6757,6734,6711,6688,6666,6643,6620,6597,6574,6550,6527,6504,6481,6458,6435,6412,6389,6366,6342,6319,6296,6273,6250,6226,6203,6180,6156,6133,6110,6086,6063,6040,6016,5993,5970,5946,5923,5899,5876,5852,5829,5805,5782,5758,5735,5711,5688,5664,5640,5617,5593,5570,5546,5522,5499,5475,5451,5427,5404,5380,5356,5332,5309,5285,5261,5237,5213,5190,5166,5142,5118,5094,5070,5046,5022,4998,4974,4950,4926,4902,4878,4854,4830,4806,4782,4758,4734,4710,4686,4662,4638,4614,4590,4565,4541,4517,4493,4469,4445,4420,4396,4372,4348,4323,4299,4275,4251,4226,4202,4178,4153,4129,4105,4080,4056,4032,4007,3983,3958,3934,3910,3885,3861,3836,3812,3787,3763,3739,3714,3690,3665,3641,3616,3591,3567,3542,3518,3493,3469,3444,3420,3395,3370,3346,3321,3296,3272,3247,3223,3198,3173,3149,3124,3099,3075,3050,3025,3000,2976,2951,2926,2901,2877,2852,2827,2802,2778,2753,2728,2703,2678,2654,2629,2604,2579,2554,2529,2505,2480,2455,2430,2405,2380,2355,2331,2306,2281,2256,2231,2206,2181,2156,2131,2106,2081,2056,2032,2007,1982,1957,1932,1907,1882,1857,1832,1807,1782,1757,1732,1707,1682,1657,1632,1607,1582,1557,1532,1507,1482,1456,1431,1406,1381,1356,1331,1306,1281,1256,1231,1206,1181,1156,1131,1106,1080,1055,1030,1005,980,955,930,905,880,855,829,804,779,754,729,704,679,654,628,603,578,553,528,503,478,453,427,402,377,352,327,302,277,251,226,201,176,151,126,101,75,50,25,0
	);

	SIGNAL sin , cos : S16;
	--SIGNAL sin , cos : S16S;

BEGIN

	sin_read: PROCESS (clk)
		--variable w_sen : U9 := 0;
	BEGIN
		IF falling_edge(clk) THEN
			sin <=  sin_rom(w);
			--sin <= to_signed(sin_rom(w),16); -- Read from ROM
			--w_sen := w;
			--while(w_sen>(sin_rom'length-1)) loop
			--	w_sen := (sin_rom'length-1) - (w_sen - (sin_rom'length-1));
			--	if (w_sen < 0) then
			--		w_sen := -w_sen;
			--	end if;
			--end loop;
			--sin <= to_signed(sin_rom(w_sen),16);
		END IF;
	END PROCESS;

	cos_read: PROCESS (clk)
		--variable w_cos : U9 := 0;
	BEGIN
		IF falling_edge(clk) THEN
			cos <=  cos_rom(w);
			--cos <=  to_signed(cos_rom(w),16); -- Read from ROM
			--w_cos := w;
			--while(w_cos>cos_rom'length-1) loop
			--	w_cos := (cos_rom'length-1) - (w_cos - (cos_rom'length-1));
			--	if (w_cos < 0) then
			--		w_cos := -w_cos;
			--	end if;
			--end loop;
			--cos <= to_signed(cos_rom(w_cos),16);
		END IF;
	END PROCESS;

	States: PROCESS(clk, reset, w)-----> FFT in behavioral style
		VARIABLE i1, i2, gcount, k1, k2   : U9 := 0;
		VARIABLE stage, dw, count, rcount  : U9 := 0;
		VARIABLE tr, ti : S16 := 0;
		--VARIABLE tr, ti : S16S := (others => '0');
		VARIABLE slv, rslv : STD_LOGIC_VECTOR(0 TO ldN-1);
	BEGIN	
		IF reset = '0' THEN  -- Asynchronous reset
			s <= start;
			fftr <= 0;
			ffti <=	0;
			--fftr <= (others => '0');
			--ffti <= (others => '0');
		ELSIF rising_edge(clk) THEN
			CASE s IS   -- Next State assignments
				WHEN start =>
					s <= load;
					count := 0;
					gcount := 0; 
					stage:= 1; 
					i1:=0; 
					i2 := N/2; 
					k1:=N;
					k2:=N/2; 
					dw := 1; 
					fft_valid <= '0';
				WHEN load =>       -- Read in all data from I/O ports
					xr(count) <= xr_in; 
					xi(count) <= xi_in;
					--xr(count) <= signed(xr_in); 
					--xi(count) <= signed(xi_in);
					count := count + 1;
					IF count = N THEN  s <= calc;
					ELSE               s <= load;
					END IF;
				WHEN calc =>          -- Do the butterfly computation
					tr := xr(i1) - xr(i2);
					xr(i1) <= xr(i1) + xr(i2);
					ti := xi(i1) - xi(i2);
					xi(i1) <= xi(i1) + xi(i2);
					xr(i2) <= (cos * tr + sin * ti)/2**14;
					xi(i2) <= (cos * ti - sin * tr)/2**14;
					--xr(i2) <= resize(shift_right((cos * tr + sin * ti),14),16);		
					--xi(i2) <= resize(shift_right((cos * ti - sin * tr),14),16);												
					s <= update;
				WHEN update =>           -- All counters and pointers
					s  <= calc; -- By default do next butterfly
					i1 := i1 + k1; -- Next butterfly in group
					i2 := i1 + k2;
					wo <= 1;
					IF i1 >= N-1 THEN -- All butterflies done in group?
						gcount := gcount + 1;
						i1 := gcount;
						i2 := i1 + k2;
						wo <= 2;
						IF gcount >= k2 THEN-- All groups done in stages?
							gcount := 0; 
							i1 := 0; 
							i2 := k2;
							dw := dw * 2;
							stage  := stage + 1;
							wo <= 3;
							IF stage > ldN THEN -- All stages done
								s <= reverse;
								count := 0;
								wo <= 4;
							ELSE -- Start new stage
								k1 := k2; k2 := k2/2;
								i1 := 0; i2 := k2;
								w<=0;wo <= 5;
							END IF;
						ELSE -- Start new group
							i1 := gcount;  i2 := i1 + k2;
							w<=w+dw;
							wo <= 6;
						END IF;
					END IF;
				WHEN reverse =>   -- Apply bitreverse
					fft_valid <= '1';
					slv := STD_LOGIC_VECTOR(to_unsigned(count, ldn));
					FOR i IN 0 TO ldn-1 LOOP
						rslv(i) := slv(ldn-i-1);
					END LOOP;
					rcount := CONV_INTEGER('0' & rslv);

					fftr <= xr(rcount);
					ffti <= xi(rcount);
					--fftr <= std_logic_vector(xr(rcount));
					--ffti <= std_logic_vector(xi(rcount));
					count := count + 1;
					IF count >= N THEN  s <= done;
					ELSE                s <= reverse;
					END IF;
				WHEN done =>      -- Output of results
					s <= start;     -- Start next cycle
			END CASE;
		END IF;
		i1_o<=i1;   -- Provide some test signals as outputs
		i2_o<=i2;
		stage_o<=stage;
		gcount_o <= gcount;
		k1_o <= k1;
		k2_o<=k2;
		w_o<=w;
		dw_o<=dw;
		rcount_o <= rcount;
	END PROCESS States;
	
	Rk: FOR k IN 0 TO 7 GENERATE -- Show first 8
		--xr_out(k) <= std_logic_vector(xr(k));        -- register values
		--xi_out(k) <= std_logic_vector(xi(k));
		xr_out(k) <= xr(k);
		xi_out(k) <= xi(k);
	END GENERATE;
	
END fpga; 
